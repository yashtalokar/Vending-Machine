interface vending_if(input logic clk);
  logic five_rup, ten_rup,reset;
  logic [3:0] item_no;
  logic product, change;
endinterface
